library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.env.finish;

ENTITY tb_cpu IS
END ENTITY;

ARCHITECTURE tb_cpu_arch OF tb_cpu IS
BEGIN
	test : PROCESS
	BEGIN
		finish;
	END PROCESS;
END ARCHITECTURE;


